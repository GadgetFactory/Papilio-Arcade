library ieee;
  use ieee.std_logic_1164.all;
  use ieee.std_logic_unsigned.all;
  use ieee.numeric_std.all;

package pkg_galaxian is
end;

package body pkg_galaxian is
end;
