library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity cart_rom is
   port(clk: in std_logic;
        d: out std_logic_vector(7 downto 0);
        a: in std_logic_vector(12 downto 0));
end cart_rom;

architecture arch of cart_rom is
   type rom_type is array (0 to 8191) of std_logic_vector(7 downto 0);
   signal rom: rom_type := (
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00");

   signal ra: std_logic_vector(12 downto 0);

begin
   process(clk)
   begin
      if (clk = '0' and clk'event) then
         ra <= a;
      end if;
   end process;

   d <= rom(to_integer(unsigned(ra)));
end arch;
